library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package instruction_buffer_type is
	constant data_size : integer := 32;  --bits wide
	constant num_of_inputs    : integer := 32; --bits wide
	constant log2_Of_num_of_inputs : integer := 5;
	type inputVectors is array(0 to num_of_inputs) of std_logic_vector (0 to data_size);
	type internalCarry is array(0 to log2_Of_num_of_inputs+1) of inputVectors;
end package instruction_buffer_type;

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.math_real.all;

use work.instruction_buffer_type.all;

entity registerFile_nbit_struct is
    -- If you cange n you must remake the decoder function
  generic(N : integer := 32);
  port(
     


    i_rd               : in std_logic_vector(0 to N);
    in_select_rs       : in std_logic_vector(0 to 5);
    in_select_rt       : in std_logic_vector(0 to 5);
    in_select_rd       : in std_logic_vector(0 to 5);
    i_WE               : in std_logic;
    i_CLK              : in std_logic;
    i_RST              : in std_logic;


    o_rt               : out std_logic_vector(0 to N);
    o_rs               : out std_logic_vector(0 to N);
    o_carry            : out std_logic

	);
	
end registerFile_nbit_struct;

architecture registerFile_nbit_struct_arch of registerFile_nbit_struct is

        signal inter_select  : std_logic_vector(0 to N);

        --G00: for i in 0 to N generate
            signal inter_carry      : inputVectors;
        --end generate;
	signal write_enable_vector : std_logic_vector(0 to N);


	component andg2
		port(
			i_A          : in std_logic;
       			i_B          : in std_logic;
       			o_F          : out std_logic
			);
	end component;
		



        component decoder5to32_flow
            port(
                i_data        : in std_logic_vector(0 to 5);     
                o_data        : in std_logic_vector(0 to 32)
                );
        end component;


        component mux_nbit_nbitto1_struct
            port(
--                G0: for i in 0 to N generate
                    in_data_0    : in inputVectors;
            
--                end generate;
            
                in_select        : in std_logic_vector(0 to 5);
                o_z              : out std_logic_vector(0 to N)


                );
        end component;


        component register_nbit_struct
            port(
                i_CLK             : in std_logic;
                i_RST             : in std_logic;
                i_WE              : in std_logic;
                i_D               : in std_logic_vector(0 to N);   
            
                o_Q               : out std_logic_vector(0 to N)
                );
        end component;

    begin

        
    -- Everything but this circuit can scale up YOU MUST REBUILD THIS TO CHANGE N
    inverter: decoder5to32_flow 
        port map(
                    i_data   => in_select_rd,
                    o_data      => inter_select     
                );



    G1: for j in 0 to N generate
            and_j: andg2
            port map(


			i_A          => inter_select(j),
       			i_B          => i_WE,
       			o_F          => write_enable_vector(j)

            );
    end generate;









    --create all of registers
    G0: for j in 0 to N generate
            register_j: register_nbit_struct
            port map(


                i_CLK             => i_CLK,
                i_RST             => i_RST,
                i_WE              => write_enable_vector(j), --only write when global write is on and this register selected 
                i_D               => i_rd,   
            
                o_Q               => inter_carry(j)

            );
    end generate;

        

    -- mux to output the rt data
    mux_rt: mux_nbit_nbitto1_struct
    port map(

            --get all the inputs from the registers
 --           G2: for i in 0 to N generate
                in_data_0    => inter_carry,
        
 --           end generate;
        
            in_select            => in_select_rt,
            o_z                  => o_rt
    );




    -- mux to output the rs data
    mux_rs: mux_nbit_nbitto1_struct
    port map(


                in_data_0    => inter_carry,
        

            in_select            => in_select_rs,
            o_z                  => o_rs
    );


        






end registerFile_nbit_struct_arch;