entity ALUcontrol is 
    port(  
        i_instructions          : in std_logic_vector(0 to 5);
        ALUctl_signal           : in std_logic_vector(0 to 4);

        ALUOpIn                 : in std_logic_vector(0 to 4)

    );

end ALUcontrol;














