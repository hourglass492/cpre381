



-- problem 4 b



entity sys2 is
    port (
        input_w     : in std_logic;
        a_data      : in std_logic_vector(0 to 7);
        b_data      : in std_logic_vector(0 to 7);
        clik        : in std_logic;
        dat_4       : out std_logic_vector(0 to 7);
        dat_4       : out std_logic_vector(0 to 3);
    );
end sys2;





